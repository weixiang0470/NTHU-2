`timescale 1ns / 1ps

module Buffer(
    input clk,
    input rst,
    input arbiter_result,
    input arbiter_done,
    output reg [7:0] response,
    output reg ready,
    output reg buf_rst
);
    // -------------------------------------------------------------------------
    // Module Declaration:
    // The Buffer module accumulates bits given by 'arbiter_result' into an
    // 8-bit 'response'. Once enough bits have been collected, 'ready' is
    // asserted to signal that the response is valid. Meanwhile, 'buf_rst'
    // can be used to reset counters and arbiters whenever a new bit is captured.
    //
    // Inputs:
    //   - clk           : clock signal for synchronous operations
    //   - rst           : active-high reset signal, clearing the module state
    //   - arbiter_result: single-bit data from race_arbiter to be stored
    //   - arbiter_done  : indicates when new arbiter_result is available
    // Outputs:
    //   - response [7:0]: the assembled bits from arbiter_result
    //   - ready         : indicates response is fully populated
    //   - buf_rst       : resets external modules while collecting bits
    // -------------------------------------------------------------------------

    // 1. Declare a register to track how many bits have been accumulated.

    // 2. Implement a synchronous block (always @(posedge clk or posedge rst)):
    //    - If rst is asserted, clear 'response', 'ready', 'buf_rst', and the counter.
    //    - Set 'ready' once the counter has reached its threshold (e.g., 7 for 8 bits).
    //    - Shift in 'arbiter_result' into 'response'.
    //    - Assert 'buf_rst' to reset external modules while a new bit is recorded.
    reg [2:0] bit_count;

    always@(posedge clk or posedge rst)begin
        if(rst) begin
            response <= 8'b0;
            ready <= 0;
            buf_rst <= 1;
            bit_count <= 0;
        end else if (arbiter_done) begin
            buf_rst <= 1;
            response <= {response[6:0], arbiter_result};
            bit_count <= bit_count + 1;
            if (bit_count == 7) begin
                ready <= 1;
                //bit_count <= 0;
            end else begin
                ready <= 0;
            end
        end else begin
            buf_rst <= 0;
        end
        
    end

endmodule