`timescale 1ns / 1ps

// module hamming_distance (
//     input [7:0] S1,  // 8-bit 输入信号 1
//     input [7:0] S2,  // 8-bit 输入信号 2
//     output reg [3:0] HD // 海明距离
// );

//     integer i;
    
//     always @(*) begin
//         HD = 0;  // 初始化海明距离
//         for (i = 0; i < 8; i = i + 1) begin
//             if (S1[i] == 1 && S2[i] == 1) begin
//                 HD = HD + 1;  // 如果同一位上 S1 和 S2 都为 1，海明距离加 1
//             end
//         end
//     end
// endmodule


module UQ_tb();

localparam real DELAY_SETS0 [0:15][0:10] = '{
    '{0.42, 0.67, 0.58, 0.88, 0.54, 0.63, 0.77, 0.45, 0.69, 0.51, 0.76},
    '{0.51, 0.81, 0.60, 0.72, 0.64, 0.85, 0.59, 0.62, 0.66, 0.79, 0.57},
    '{0.79, 0.66, 0.61, 0.55, 0.56, 0.69, 0.51, 0.68, 0.70, 0.63, 0.73},
    '{0.53, 0.58, 0.63, 0.55, 0.52, 0.77, 0.69, 0.61, 0.79, 0.62, 0.78},
    '{0.66, 0.70, 0.81, 0.60, 0.52, 0.68, 0.64, 0.74, 0.72, 0.58, 0.55},
    '{0.72, 0.56, 0.54, 0.68, 0.62, 0.80, 0.51, 0.75, 0.82, 0.74, 0.56},
    '{0.59, 0.53, 0.70, 0.71, 0.64, 0.79, 0.65, 0.73, 0.57, 0.67, 0.69},
    '{0.61, 0.66, 0.67, 0.78, 0.80, 0.52, 0.54, 0.65, 0.66, 0.72, 0.74},
    '{0.75, 0.62, 0.67, 0.56, 0.58, 0.68, 0.61, 0.73, 0.78, 0.53, 0.67},
    '{0.87, 0.62, 0.39, 0.92, 0.73, 0.51, 0.64, 0.71, 0.56, 0.43, 0.76},
    '{0.64, 0.60, 0.77, 0.75, 0.69, 0.72, 0.62, 0.57, 0.65, 0.61, 0.58},
    '{0.55, 0.72, 0.69, 0.53, 0.57, 0.78, 0.80, 0.71, 0.76, 0.59, 0.64},
    '{0.69, 0.58, 0.76, 0.75, 0.63, 0.65, 0.59, 0.74, 0.67, 0.70, 0.66},
    '{0.60, 0.66, 0.62, 0.55, 0.80, 0.68, 0.73, 0.72, 0.67, 0.78, 0.69},
    '{0.70, 0.56, 0.54, 0.58, 0.74, 0.80, 0.52, 0.69, 0.62, 0.66, 0.60},
    '{0.74, 0.67, 0.64, 0.62, 0.59, 0.69, 0.76, 0.55, 0.60, 0.67, 0.73}
};

localparam real DELAY_SETS1 [0:15][0:10] = '{
    '{0.49, 0.62, 0.69, 0.71, 0.55, 0.67, 0.53, 0.61, 0.73, 0.64, 0.79},
    '{0.55, 0.77, 0.68, 0.34, 0.82, 0.58, 0.67, 0.64, 0.79, 0.92, 0.69},
    '{0.50, 0.74, 0.60, 0.80, 0.68, 0.55, 0.58, 0.67, 0.79, 0.62, 0.70},
    '{0.65, 0.54, 0.69, 0.72, 0.63, 0.67, 0.55, 0.70, 0.62, 0.77, 0.56},
    '{0.66, 0.53, 0.60, 0.68, 0.76, 0.80, 0.72, 0.64, 0.57, 0.59, 0.75},
    '{0.57, 0.67, 0.72, 0.61, 0.64, 0.66, 0.69, 0.53, 0.55, 0.58, 0.78},
    '{0.68, 0.71, 0.62, 0.56, 0.67, 0.69, 0.75, 0.71, 0.55, 0.74, 0.77},
    '{0.65, 0.74, 0.59, 0.56, 0.63, 0.62, 0.68, 0.60, 0.69, 0.74, 0.73},
    '{0.56, 0.79, 0.64, 0.66, 0.61, 0.68, 0.67, 0.61, 0.55, 0.58, 0.69},
    '{0.57, 0.64, 0.70, 0.65, 0.60, 0.67, 0.58, 0.61, 0.75, 0.78, 0.72},
    '{0.63, 0.55, 0.80, 0.59, 0.61, 0.70, 0.52, 0.58, 0.63, 0.74, 0.67},
    '{0.59, 0.73, 0.56, 0.72, 0.61, 0.79, 0.68, 0.62, 0.56, 0.69, 0.75},
    '{0.68, 0.54, 0.72, 0.67, 0.79, 0.59, 0.60, 0.63, 0.66, 0.55, 0.74},
    '{0.64, 0.72, 0.70, 0.59, 0.62, 0.69, 0.74, 0.61, 0.56, 0.72, 0.55},
    '{0.56, 0.60, 0.68, 0.57, 0.63, 0.64, 0.75, 0.77, 0.73, 0.56, 0.72},
    '{0.74, 0.58, 0.61, 0.69, 0.63, 0.57, 0.68, 0.74, 0.70, 0.79, 0.60}
};

localparam real DELAY_SETS2 [0:15][0:10] = '{
    '{0.73, 0.72, 0.60, 0.68, 0.55, 0.76, 0.77, 0.62, 0.64, 0.69, 0.72},
    '{0.65, 0.71, 0.62, 0.60, 0.78, 0.64, 0.58, 0.66, 0.75, 0.68, 0.80},
    '{0.62, 0.72, 0.66, 0.63, 0.71, 0.70, 0.69, 0.65, 0.55, 0.57, 0.66},
    '{0.54, 0.61, 0.60, 0.75, 0.74, 0.56, 0.59, 0.67, 0.68, 0.62, 0.65},
    '{0.61, 0.57, 0.64, 0.75, 0.72, 0.78, 0.59, 0.63, 0.56, 0.70, 0.71},
    '{0.75, 0.65, 0.60, 0.64, 0.56, 0.62, 0.59, 0.57, 0.74, 0.69, 0.68},
    '{0.34, 0.78, 0.56, 0.49, 0.71, 0.58, 0.65, 0.72, 0.81, 0.66, 0.80},
    '{0.60, 0.59, 0.71, 0.56, 0.72, 0.64, 0.75, 0.66, 0.70, 0.73, 0.71},
    '{0.62, 0.55, 0.70, 0.64, 0.61, 0.68, 0.72, 0.78, 0.75, 0.68, 0.61},
    '{0.74, 0.67, 0.66, 0.59, 0.71, 0.75, 0.79, 0.63, 0.77, 0.66, 0.60},
    '{0.62, 0.75, 0.64, 0.59, 0.80, 0.71, 0.68, 0.60, 0.72, 0.73, 0.64},
    '{0.67, 0.56, 0.70, 0.63, 0.74, 0.60, 0.65, 0.72, 0.69, 0.61, 0.63},
    '{0.75, 0.61, 0.72, 0.67, 0.59, 0.67, 0.62, 0.70, 0.65, 0.75, 0.71},
    '{0.63, 0.59, 0.65, 0.72, 0.70, 0.62, 0.68, 0.61, 0.60, 0.58, 0.63},
    '{0.74, 0.68, 0.56, 0.65, 0.72, 0.60, 0.77, 0.55, 0.67, 0.63, 0.72},
    '{0.61, 0.65, 0.74, 0.62, 0.75, 0.59, 0.68, 0.60, 0.69, 0.77, 0.63}
};

localparam real DELAY_SETS3 [0:15][0:10] = '{
    '{0.52, 0.67, 0.72, 0.74, 0.56, 0.64, 0.58, 0.79, 0.75, 0.62, 0.61},
    '{0.69, 0.65, 0.59, 0.80, 0.92, 0.49, 0.77, 0.51, 0.75, 0.50, 0.68},
    '{0.71, 0.66, 0.65, 0.57, 0.75, 0.59, 0.63, 0.77, 0.58, 0.73, 0.69},
    '{0.59, 0.66, 0.54, 0.72, 0.70, 0.63, 0.61, 0.68, 0.77, 0.74, 0.55},
    '{0.67, 0.59, 0.74, 0.62, 0.75, 0.80, 0.68, 0.71, 0.64, 0.55, 0.56},
    '{0.63, 0.76, 0.59, 0.67, 0.60, 0.68, 0.70, 0.57, 0.74, 0.76, 0.80},
    '{0.62, 0.71, 0.65, 0.66, 0.75, 0.80, 0.66, 0.59, 0.58, 0.63, 0.65},
    '{0.77, 0.75, 0.69, 0.74, 0.70, 0.66, 0.61, 0.62, 0.78, 0.61, 0.59},
    '{0.55, 0.64, 0.79, 0.68, 0.60, 0.62, 0.73, 0.77, 0.68, 0.72, 0.71},
    '{0.60, 0.69, 0.77, 0.64, 0.74, 0.67, 0.76, 0.65, 0.72, 0.75, 0.79},
    '{0.70, 0.62, 0.55, 0.71, 0.73, 0.79, 0.58, 0.78, 0.69, 0.60, 0.77},
    '{0.64, 0.61, 0.66, 0.56, 0.61, 0.78, 0.70, 0.58, 0.72, 0.65, 0.65},
    '{0.55, 0.76, 0.60, 0.65, 0.79, 0.67, 0.58, 0.74, 0.69, 0.74, 0.72},
    '{0.66, 0.73, 0.70, 0.72, 0.64, 0.55, 0.67, 0.62, 0.61, 0.69, 0.59},
    '{0.75, 0.67, 0.74, 0.63, 0.72, 0.71, 0.55, 0.65, 0.63, 0.59, 0.75},
    '{0.60, 0.61, 0.58, 0.75, 0.69, 0.66, 0.61, 0.72, 0.64, 0.75, 0.70}
};

localparam real DELAY_SETS4 [0:15][0:10] = '{
    '{0.64, 0.60, 0.67, 0.72, 0.56, 0.69, 0.62, 0.78, 0.73, 0.66, 0.58},
    '{0.68, 0.71, 0.66, 0.75, 0.63, 0.64, 0.58, 0.77, 0.79, 0.66, 0.65},
    '{0.67, 0.75, 0.58, 0.60, 0.70, 0.72, 0.65, 0.68, 0.66, 0.75, 0.69},
    '{0.62, 0.61, 0.78, 0.64, 0.55, 0.59, 0.63, 0.67, 0.72, 0.56, 0.79},
    '{0.77, 0.60, 0.56, 0.72, 0.67, 0.73, 0.75, 0.62, 0.68, 0.77, 0.61},
    '{0.68, 0.61, 0.59, 0.64, 0.76, 0.73, 0.60, 0.79, 0.66, 0.65, 0.55},
    '{0.70, 0.77, 0.65, 0.66, 0.60, 0.71, 0.74, 0.69, 0.72, 0.75, 0.63},
    '{0.55, 0.67, 0.62, 0.71, 0.64, 0.63, 0.67, 0.65, 0.70, 0.66, 0.75},
    '{0.79, 0.64, 0.67, 0.75, 0.61, 0.74, 0.78, 0.72, 0.62, 0.65, 0.68},
    '{0.68, 0.60, 0.72, 0.67, 0.63, 0.64, 0.78, 0.66, 0.75, 0.55, 0.73},
    '{0.62, 0.55, 0.63, 0.66, 0.79, 0.61, 0.60, 0.67, 0.75, 0.64, 0.72},
    '{0.61, 0.72, 0.70, 0.59, 0.75, 0.68, 0.66, 0.73, 0.60, 0.68, 0.65},
    '{0.79, 0.55, 0.64, 0.72, 0.66, 0.58, 0.77, 0.63, 0.75, 0.68, 0.74},
    '{0.60, 0.59, 0.73, 0.52, 0.61, 0.67, 0.80, 0.79, 0.68, 0.76, 0.71},
    '{0.60, 0.72, 0.68, 0.66, 0.73, 0.75, 0.70, 0.56, 0.74, 0.61, 0.67},
    '{0.69, 0.64, 0.60, 0.66, 0.71, 0.74, 0.55, 0.61, 0.72, 0.67, 0.58}
};

localparam real DELAY_SETS5 [0:15][0:10] = '{
    '{0.66, 0.68, 0.60, 0.73, 0.71, 0.77, 0.56, 0.63, 0.58, 0.62, 0.67},
    '{0.61, 0.72, 0.67, 0.66, 0.75, 0.73, 0.79, 0.70, 0.63, 0.64, 0.55},
    '{0.81, 0.62, 0.65, 0.72, 0.55, 0.61, 0.63, 0.74, 0.77, 0.56, 0.78},
    '{0.74, 0.77, 0.62, 0.60, 0.69, 0.72, 0.73, 0.61, 0.67, 0.75, 0.79},
    '{0.70, 0.61, 0.63, 0.65, 0.75, 0.67, 0.61, 0.77, 0.72, 0.65, 0.79},
    '{0.64, 0.74, 0.78, 0.59, 0.70, 0.76, 0.73, 0.75, 0.62, 0.79, 0.67},
    '{0.59, 0.66, 0.75, 0.62, 0.68, 0.73, 0.55, 0.77, 0.74, 0.64, 0.68},
    '{0.65, 0.68, 0.60, 0.66, 0.72, 0.63, 0.71, 0.65, 0.66, 0.78, 0.56},
    '{0.75, 0.67, 0.69, 0.61, 0.79, 0.60, 0.72, 0.74, 0.66, 0.61, 0.62},
    '{0.74, 0.75, 0.63, 0.70, 0.72, 0.68, 0.60, 0.66, 0.75, 0.69, 0.67},
    '{0.60, 0.66, 0.62, 0.69, 0.68, 0.72, 0.77, 0.75, 0.59, 0.64, 0.63},
    '{0.64, 0.68, 0.71, 0.73, 0.75, 0.78, 0.52, 0.53, 0.69, 0.56, 0.85},
    '{0.69, 0.65, 0.76, 0.74, 0.67, 0.62, 0.61, 0.70, 0.75, 0.64, 0.58},
    '{0.61, 0.78, 0.69, 0.63, 0.66, 0.74, 0.60, 0.61, 0.55, 0.64, 0.72},
    '{0.63, 0.75, 0.71, 0.62, 0.59, 0.75, 0.67, 0.71, 0.74, 0.79, 0.69},
    '{0.65, 0.62, 0.76, 0.69, 0.74, 0.67, 0.60, 0.77, 0.59, 0.70, 0.67}
};

localparam real DELAY_SETS6 [0:15][0:10] = '{
    '{0.74, 0.79, 0.72, 0.67, 0.73, 0.60, 0.61, 0.68, 0.66, 0.75, 0.78},
    '{0.56, 0.67, 0.70, 0.72, 0.75, 0.60, 0.62, 0.76, 0.63, 0.75, 0.74},
    '{0.64, 0.61, 0.62, 0.67, 0.66, 0.60, 0.65, 0.78, 0.75, 0.69, 0.68},
    '{0.63, 0.71, 0.85, 0.47, 0.59, 0.77, 0.55, 0.62, 0.66, 0.64, 0.48},
    '{0.75, 0.69, 0.72, 0.59, 0.68, 0.61, 0.60, 0.64, 0.73, 0.72, 0.77},
    '{0.69, 0.65, 0.66, 0.61, 0.75, 0.70, 0.67, 0.64, 0.63, 0.71, 0.72},
    '{0.67, 0.79, 0.65, 0.72, 0.74, 0.75, 0.67, 0.66, 0.76, 0.60, 0.67},
    '{0.72, 0.70, 0.73, 0.61, 0.63, 0.67, 0.69, 0.75, 0.61, 0.59, 0.74},
    '{0.55, 0.67, 0.69, 0.54, 0.73, 0.66, 0.70, 0.63, 0.79, 0.59, 0.57},
    '{0.75, 0.72, 0.67, 0.65, 0.66, 0.60, 0.61, 0.78, 0.71, 0.74, 0.75},
    '{0.60, 0.64, 0.62, 0.77, 0.71, 0.78, 0.69, 0.73, 0.62, 0.59, 0.64},
    '{0.79, 0.70, 0.67, 0.74, 0.62, 0.65, 0.61, 0.73, 0.64, 0.69, 0.61},
    '{0.75, 0.63, 0.67, 0.66, 0.60, 0.74, 0.69, 0.75, 0.61, 0.72, 0.64},
    '{0.63, 0.62, 0.65, 0.66, 0.67, 0.75, 0.70, 0.67, 0.64, 0.75, 0.70},
    '{0.75, 0.66, 0.68, 0.74, 0.62, 0.75, 0.68, 0.63, 0.72, 0.66, 0.74},
    '{0.67, 0.76, 0.72, 0.60, 0.68, 0.71, 0.73, 0.75, 0.78, 0.66, 0.65}
};

localparam real DELAY_SETS7 [0:15][0:10] = '{
    '{0.62, 0.73, 0.66, 0.74, 0.60, 0.68, 0.70, 0.75, 0.77, 0.64, 0.72},
    '{0.69, 0.68, 0.63, 0.75, 0.74, 0.66, 0.72, 0.67, 0.71, 0.73, 0.70},
    '{0.66, 0.77, 0.62, 0.72, 0.65, 0.70, 0.74, 0.61, 0.69, 0.75, 0.67},
    '{0.75, 0.64, 0.68, 0.72, 0.70, 0.63, 0.69, 0.67, 0.74, 0.71, 0.78},
    '{0.67, 0.62, 0.60, 0.75, 0.64, 0.72, 0.78, 0.71, 0.73, 0.75, 0.68},
    '{0.66, 0.70, 0.67, 0.63, 0.74, 0.79, 0.75, 0.71, 0.72, 0.68, 0.76},
    '{0.74, 0.65, 0.69, 0.72, 0.70, 0.68, 0.63, 0.75, 0.64, 0.77, 0.71},
    '{0.77, 0.69, 0.71, 0.75, 0.66, 0.72, 0.79, 0.70, 0.60, 0.65, 0.74},
    '{0.61, 0.75, 0.74, 0.68, 0.66, 0.72, 0.63, 0.77, 0.67, 0.69, 0.64},
    '{0.63, 0.61, 0.75, 0.55, 0.80, 0.59, 0.71, 0.60, 0.72, 0.54, 0.79},
    '{0.70, 0.64, 0.66, 0.72, 0.61, 0.69, 0.74, 0.65, 0.68, 0.75, 0.62},
    '{0.72, 0.71, 0.65, 0.74, 0.70, 0.73, 0.67, 0.79, 0.76, 0.68, 0.61},
    '{0.63, 0.71, 0.69, 0.66, 0.70, 0.75, 0.74, 0.66, 0.72, 0.67, 0.73},
    '{0.75, 0.74, 0.63, 0.61, 0.77, 0.72, 0.78, 0.66, 0.73, 0.68, 0.65},
    '{0.74, 0.63, 0.69, 0.77, 0.62, 0.72, 0.70, 0.65, 0.73, 0.68, 0.75},
    '{0.76, 0.67, 0.72, 0.61, 0.70, 0.65, 0.67, 0.63, 0.72, 0.69, 0.71}
};

localparam real DELAY_SETS8 [0:15][0:10] = '{
    '{0.70, 0.61, 0.75, 0.72, 0.67, 0.63, 0.79, 0.74, 0.71, 0.77, 0.62},
    '{0.73, 0.75, 0.66, 0.71, 0.70, 0.72, 0.63, 0.64, 0.68, 0.79, 0.67},
    '{0.61, 0.65, 0.71, 0.74, 0.69, 0.72, 0.63, 0.79, 0.75, 0.77, 0.64},
    '{0.72, 0.68, 0.60, 0.75, 0.66, 0.70, 0.77, 0.71, 0.79, 0.68, 0.67},
    '{0.66, 0.65, 0.62, 0.68, 0.75, 0.61, 0.70, 0.63, 0.79, 0.72, 0.64},
    '{0.63, 0.74, 0.67, 0.79, 0.61, 0.72, 0.74, 0.71, 0.63, 0.70, 0.75},
    '{0.66, 0.65, 0.74, 0.72, 0.67, 0.61, 0.71, 0.70, 0.75, 0.64, 0.76},
    '{0.75, 0.72, 0.67, 0.62, 0.55, 0.66, 0.70, 0.68, 0.64, 0.59, 0.73},
    '{0.71, 0.75, 0.63, 0.68, 0.67, 0.62, 0.74, 0.77, 0.70, 0.79, 0.66},
    '{0.77, 0.64, 0.69, 0.75, 0.66, 0.73, 0.74, 0.62, 0.79, 0.65, 0.71},
    '{0.65, 0.72, 0.75, 0.79, 0.61, 0.66, 0.63, 0.70, 0.69, 0.74, 0.60},
    '{0.75, 0.70, 0.74, 0.64, 0.72, 0.67, 0.79, 0.73, 0.71, 0.65, 0.63},
    '{0.70, 0.63, 0.75, 0.67, 0.72, 0.60, 0.74, 0.66, 0.68, 0.69, 0.71},
    '{0.69, 0.66, 0.75, 0.63, 0.60, 0.72, 0.79, 0.64, 0.68, 0.71, 0.65},
    '{0.62, 0.70, 0.77, 0.74, 0.63, 0.75, 0.71, 0.78, 0.65, 0.68, 0.72},
    '{0.74, 0.76, 0.69, 0.70, 0.67, 0.72, 0.63, 0.75, 0.79, 0.77, 0.66}
};

localparam real DELAY_SETS9 [0:15][0:10] = '{
    '{0.70, 0.75, 0.74, 0.65, 0.69, 0.63, 0.62, 0.77, 0.76, 0.61, 0.64},
    '{0.67, 0.61, 0.68, 0.71, 0.75, 0.74, 0.64, 0.70, 0.79, 0.76, 0.75},
    '{0.73, 0.76, 0.77, 0.74, 0.72, 0.75, 0.63, 0.72, 0.70, 0.78, 0.64},
    '{0.75, 0.71, 0.79, 0.74, 0.68, 0.72, 0.60, 0.77, 0.65, 0.67, 0.69},
    '{0.73, 0.74, 0.71, 0.69, 0.70, 0.75, 0.76, 0.62, 0.79, 0.64, 0.66},
    '{0.74, 0.68, 0.77, 0.65, 0.71, 0.62, 0.78, 0.75, 0.67, 0.74, 0.73},
    '{0.61, 0.76, 0.72, 0.69, 0.70, 0.64, 0.78, 0.75, 0.61, 0.73, 0.77},
    '{0.67, 0.75, 0.64, 0.73, 0.70, 0.76, 0.75, 0.78, 0.66, 0.72, 0.74},
    '{0.71, 0.75, 0.68, 0.63, 0.79, 0.72, 0.70, 0.69, 0.76, 0.64, 0.75},
    '{0.60, 0.65, 0.66, 0.75, 0.69, 0.74, 0.78, 0.62, 0.68, 0.76, 0.71},
    '{0.78, 0.74, 0.69, 0.67, 0.61, 0.67, 0.75, 0.72, 0.62, 0.59, 0.61},
    '{0.71, 0.75, 0.64, 0.62, 0.66, 0.60, 0.57, 0.70, 0.76, 0.64, 0.68},
    '{0.75, 0.68, 0.77, 0.66, 0.72, 0.60, 0.70, 0.75, 0.67, 0.79, 0.62},
    '{0.79, 0.74, 0.73, 0.75, 0.71, 0.64, 0.69, 0.68, 0.60, 0.67, 0.75},
    '{0.70, 0.71, 0.75, 0.72, 0.69, 0.76, 0.61, 0.64, 0.79, 0.62, 0.70},
    '{0.75, 0.74, 0.77, 0.71, 0.70, 0.78, 0.69, 0.67, 0.63, 0.62, 0.75}
};

    parameter WIDTH = 3;
    
    reg clk, en, sys_rst_pos;
    reg [7:0] chall_in;
    wire [9:0][7:0] response ;
    wire [9:0]ready ;

    // Instantiate the Top module
    Top #(.DELAY_SETS(DELAY_SETS0), .WIDTH(WIDTH)) uut0 (
        .clk(clk),
        .en(en),
        .sys_rst_pos(sys_rst_pos),
        .chall_in(chall_in),
        .response(response[0]),
        .ready(ready[0])
    );
    Top #(.DELAY_SETS(DELAY_SETS1), .WIDTH(WIDTH)) uut1 (
        .clk(clk),
        .en(en),
        .sys_rst_pos(sys_rst_pos),
        .chall_in(chall_in),
        .response(response[1]),
        .ready(ready[1])
    );
    Top #(.DELAY_SETS(DELAY_SETS2), .WIDTH(WIDTH)) uut2 (
        .clk(clk),
        .en(en),
        .sys_rst_pos(sys_rst_pos),
        .chall_in(chall_in),
        .response(response[2]),
        .ready(ready[2])
    );
    Top #(.DELAY_SETS(DELAY_SETS3), .WIDTH(WIDTH)) uut3 (
        .clk(clk),
        .en(en),
        .sys_rst_pos(sys_rst_pos),
        .chall_in(chall_in),
        .response(response[3]),
        .ready(ready[3])
    );
    Top #(.DELAY_SETS(DELAY_SETS4), .WIDTH(WIDTH)) uut4 (
        .clk(clk),
        .en(en),
        .sys_rst_pos(sys_rst_pos),
        .chall_in(chall_in),
        .response(response[4]),
        .ready(ready[4])
    );
    Top #(.DELAY_SETS(DELAY_SETS5), .WIDTH(WIDTH)) uut5 (
        .clk(clk),
        .en(en),
        .sys_rst_pos(sys_rst_pos),
        .chall_in(chall_in),
        .response(response[5]),
        .ready(ready[5])
    );
    Top #(.DELAY_SETS(DELAY_SETS6), .WIDTH(WIDTH)) uut6 (
        .clk(clk),
        .en(en),
        .sys_rst_pos(sys_rst_pos),
        .chall_in(chall_in),
        .response(response[6]),
        .ready(ready[6])
    );
    Top #(.DELAY_SETS(DELAY_SETS7), .WIDTH(WIDTH)) uut7 (
        .clk(clk),
        .en(en),
        .sys_rst_pos(sys_rst_pos),
        .chall_in(chall_in),
        .response(response[7]),
        .ready(ready[7])
    );
    Top #(.DELAY_SETS(DELAY_SETS8), .WIDTH(WIDTH)) uut8 (
        .clk(clk),
        .en(en),
        .sys_rst_pos(sys_rst_pos),
        .chall_in(chall_in),
        .response(response[8]),
        .ready(ready[8])
    );
    Top #(.DELAY_SETS(DELAY_SETS9), .WIDTH(WIDTH)) uut9 (
        .clk(clk),
        .en(en),
        .sys_rst_pos(sys_rst_pos),
        .chall_in(chall_in),
        .response(response[9]),
        .ready(ready[9])
    );



    always #5 clk = ~clk;

    initial begin
        $fsdbDumpfile("UQ_tb.fsdb");
        $fsdbDumpvars(0, UQ_tb);
    end

                        

    integer hd,total_hd;
    real UQ;
    integer i, j,b;
    reg [9:0] all_ready;
    reg [9:0][7:0] all_response;
    always @(posedge ready[0])begin
        if(ready[0]) begin
            all_ready[0] = 1;
            all_response[0]=response[0];
        end
    end
    always @(posedge ready[1])begin
        if(ready[1]) begin
            all_ready[1] = 1;
            all_response[1]=response[1];
        end
    end
    always @(  posedge ready[2] ) begin
        if(ready[2]) begin
            all_ready[2] = 1;
            all_response[2]=response[2];
            // $display("Response 2 = %h",response[2]);
        end
    end
    always @(  posedge ready[3] ) begin
        if(ready[3]) begin
            all_ready[3] = 1;
            all_response[3]=response[3];
        end
    end
    always @(  posedge ready[4] ) begin
        if(ready[4]) begin
            all_ready[4] = 1;
            all_response[4]=response[4];
        end
    end
    always @(  posedge ready[5] ) begin
        if(ready[5]) begin
            all_ready[5] = 1;
            all_response[5]=response[5];
        end
    end
    always @(  posedge ready[6] ) begin
        if(ready[6]) begin
            all_ready[6] = 1;
            all_response[6]=response[6];
        end
    end
    always @(  posedge ready[7] ) begin
        if(ready[7]) begin
            all_ready[7] = 1;
            all_response[7]=response[7];
        end
    end
    always @(  posedge ready[8] ) begin
        if(ready[8]) begin
            all_ready[8] = 1;
            all_response[8]=response[8];
        end
    end
    always @(  posedge ready[9] ) begin
        if(ready[9]) begin
            all_ready[9] = 1;
            all_response[9]=response[9];
        end
    end

    always @(*) begin
        if (all_ready == 10'b1111111111) begin
            $display("CHIP 0 : at time %t, chall_in = %h, response = %h, ready = %b", $time, chall_in, all_response[0], all_ready[0]);
            $display("CHIP 1 : at time %t, chall_in = %h, response = %h, ready = %b", $time, chall_in, all_response[1], all_ready[1]);
            $display("CHIP 2 : at time %t, chall_in = %h, response = %h, ready = %b", $time, chall_in, all_response[2], all_ready[2]);
            $display("CHIP 3 : at time %t, chall_in = %h, response = %h, ready = %b", $time, chall_in, all_response[3], all_ready[3]);
            $display("CHIP 4 : at time %t, chall_in = %h, response = %h, ready = %b", $time, chall_in, all_response[4], all_ready[4]);
            $display("CHIP 5 : at time %t, chall_in = %h, response = %h, ready = %b", $time, chall_in, all_response[5], all_ready[5]);
            $display("CHIP 6 : at time %t, chall_in = %h, response = %h, ready = %b", $time, chall_in, all_response[6], all_ready[6]);
            $display("CHIP 7 : at time %t, chall_in = %h, response = %h, ready = %b", $time, chall_in, all_response[7], all_ready[7]);
            $display("CHIP 8 : at time %t, chall_in = %h, response = %h, ready = %b", $time, chall_in, all_response[8], all_ready[8]);
            $display("CHIP 9 : at time %t, chall_in = %h, response = %h, ready = %b", $time, chall_in, all_response[9], all_ready[9]);
            UQ = 0;
            total_hd=0;
            for (i=0;i<10;i=i+1)begin
                for(j=i+1;j<10;j=j+1)begin
                    hd = 0;
                    for (b = 0; b<9;b=b+1)begin
                        if(all_response[i][b] != all_response[j][b])begin
                            hd = hd+1;
                        end
                    end
                    // $display("hd = %0d",hd);
                    total_hd = total_hd + hd;
                    // $display("total_hd = %0.3f hd = %0d",total_hd,hd);
                end

            end
            UQ = (2.0/(10.0*9.0))*(total_hd / 8.0);
            $display("UQ = %0.2f",UQ);
            all_ready<=0;
        end
    end

    initial begin
        clk = 0;
        // first challenge
        $display("First challenge");

        en = 0;
        sys_rst_pos = 1;
        chall_in = 8'h01;
        #10
        sys_rst_pos = 0;
        #10
        en = 1;
        #2000

        // second challenge
        $display("Second challenge");
        en = 0;
        sys_rst_pos = 1;
        chall_in = 8'hc1;
        #10
        sys_rst_pos = 0;
        #10
        en = 1;
        #2000
        
        // third challenge
        $display("Third challenge");
        en = 0;
        sys_rst_pos = 1;
        chall_in = 8'h2c;
        #10
        sys_rst_pos = 0;
        #10
        en = 1;
        #2000
        
        // fourth challenge
        $display("Fourth challenge");
        en = 0;
        sys_rst_pos = 1;
        chall_in = 8'h01;
        #10
        sys_rst_pos = 0;
        #10
        en = 1;
        #2000

        $finish;
    end


endmodule